module nand2(x, y, s);
  input x, y;
  output s;
  
  assign s = ~(x & y);
endmodule
