module hadd(x, y, s, c);
  input x, y;
  output s, c;
  
  assign s = a ^ b;
  assign c = a & b;
endmodule